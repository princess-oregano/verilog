`ifndef OPCODE
`define OPCODE

parameter [3:0] ADD = 'd1;
parameter [3:0] SUB = 'd2;
parameter [3:0] SLL = 'd3;
parameter [3:0] SLT = 'd4;
parameter [3:0] SLTU= 'd5;
parameter [3:0] XOR = 'd6;
parameter [3:0] SRL = 'd7;
parameter [3:0] SRA = 'd8;
parameter [3:0] OR  = 'd9;
parameter [3:0] AND = 'd10;

`endif

`ifndef CMP
`define CMP

`define CMPOP_WIDTH 3
`define CMP_X       `CMPOP_WIDTH'dX
`define CMP_BEQ     `CMPOP_WIDTH'd0
`define CMP_BNE     `CMPOP_WIDTH'd1
`define CMP_BLT     `CMPOP_WIDTH'd2
`define CMP_BGE     `CMPOP_WIDTH'd3
`define CMP_BLTU    `CMPOP_WIDTH'd4
`define CMP_BGEU    `CMPOP_WIDTH'd5

`endif // CMP


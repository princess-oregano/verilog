`CASE_OP("LUI",   17'b???????_???_0110111, `ALU_X,    `ALUSEL1_X,    `ALUSEL2_X,    `WBSEL_UIMM,   1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("AUIPC", 17'b???????_???_0010111, `ALU_ADD,  `ALUSEL1_UIMM, `ALUSEL2_PC,   `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)

`CASE_OP("JAL",   17'b???????_???_1101111, `ALU_ADD,  `ALUSEL1_JIMM, `ALUSEL2_PC,   `WBSEL_PCNEXT, 1'b1, `CMP_X,    1'b0, 1'b1, 1'b0, 4'b0000)
`CASE_OP("JALR",  17'b???????_000_1100111, `ALU_ADD,  `ALUSEL1_SRC1, `ALUSEL2_IIMM, `WBSEL_PCNEXT, 1'b1, `CMP_X,    1'b0, 1'b1, 1'b0, 4'b0000)

`CASE_OP("BEQ",   17'b???????_000_1100011, `ALU_ADD,  `ALUSEL1_BIMM, `ALUSEL2_PC,   `WBSEL_X,      1'b0, `CMP_BEQ,  1'b1, 1'b0, 1'b0, 4'b0000)
`CASE_OP("BNE",   17'b???????_001_1100011, `ALU_ADD,  `ALUSEL1_BIMM, `ALUSEL2_PC,   `WBSEL_X,      1'b0, `CMP_BNE,  1'b1, 1'b0, 1'b0, 4'b0000)
`CASE_OP("BLT",   17'b???????_100_1100011, `ALU_ADD,  `ALUSEL1_BIMM, `ALUSEL2_PC,   `WBSEL_X,      1'b0, `CMP_BLT,  1'b1, 1'b0, 1'b0, 4'b0000)
`CASE_OP("BGE",   17'b???????_101_1100011, `ALU_ADD,  `ALUSEL1_BIMM, `ALUSEL2_PC,   `WBSEL_X,      1'b0, `CMP_BGE,  1'b1, 1'b0, 1'b0, 4'b0000)
`CASE_OP("BLTU",  17'b???????_110_1100011, `ALU_ADD,  `ALUSEL1_BIMM, `ALUSEL2_PC,   `WBSEL_X,      1'b0, `CMP_BLTU, 1'b1, 1'b0, 1'b0, 4'b0000)
`CASE_OP("BGEU",  17'b???????_111_1100011, `ALU_ADD,  `ALUSEL1_BIMM, `ALUSEL2_PC,   `WBSEL_X,      1'b0, `CMP_BGEU, 1'b1, 1'b0, 1'b0, 4'b0000)

`CASE_OP("LB",    17'b???????_000_0000011, `ALU_ADD,  `ALUSEL1_SRC1, `ALUSEL2_IIMM, `WBSEL_LSU,    1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("LH",    17'b???????_001_0000011, `ALU_ADD,  `ALUSEL1_SRC1, `ALUSEL2_IIMM, `WBSEL_LSU,    1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("LW",    17'b???????_010_0000011, `ALU_ADD,  `ALUSEL1_SRC1, `ALUSEL2_IIMM, `WBSEL_LSU,    1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("LBU",   17'b???????_100_0000011, `ALU_ADD,  `ALUSEL1_SRC1, `ALUSEL2_IIMM, `WBSEL_LSU,    1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("LHU",   17'b???????_101_0000011, `ALU_ADD,  `ALUSEL1_SRC1, `ALUSEL2_IIMM, `WBSEL_LSU,    1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)

`CASE_OP("SB",    17'b???????_000_0100011, `ALU_ADD,  `ALUSEL1_SRC1, `ALUSEL2_SIMM, `WBSEL_X,      1'b0, `CMP_X,    1'b0, 1'b0, 1'b1, 4'b1111)
`CASE_OP("SH",    17'b???????_001_0100011, `ALU_ADD,  `ALUSEL1_SRC1, `ALUSEL2_SIMM, `WBSEL_X,      1'b0, `CMP_X,    1'b0, 1'b0, 1'b1, 4'b1111)
`CASE_OP("SW",    17'b???????_010_0100011, `ALU_ADD,  `ALUSEL1_SRC1, `ALUSEL2_SIMM, `WBSEL_X,      1'b0, `CMP_X,    1'b0, 1'b0, 1'b1, 4'b1111)

`CASE_OP("ADDI",  17'b???????_000_0010011, `ALU_ADD,  `ALUSEL1_SRC1, `ALUSEL2_IIMM, `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("SLTI",  17'b???????_010_0010011, `ALU_SLT,  `ALUSEL1_SRC1, `ALUSEL2_IIMM, `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("SLTIU", 17'b???????_011_0010011, `ALU_SLTU, `ALUSEL1_SRC1, `ALUSEL2_IIMM, `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("XORI",  17'b???????_100_0010011, `ALU_XOR,  `ALUSEL1_SRC1, `ALUSEL2_IIMM, `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("ORI",   17'b???????_110_0010011, `ALU_OR,   `ALUSEL1_SRC1, `ALUSEL2_IIMM, `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("ANDI",  17'b???????_111_0010011, `ALU_AND,  `ALUSEL1_SRC1, `ALUSEL2_IIMM, `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("SLLI",  17'b0000000_001_0010011, `ALU_AND,  `ALUSEL1_SRC1, `ALUSEL2_IIMM, `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("SLRI",  17'b0000000_101_0010011, `ALU_AND,  `ALUSEL1_SRC1, `ALUSEL2_IIMM, `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("SRAI",  17'b0100000_101_0010011, `ALU_AND,  `ALUSEL1_SRC1, `ALUSEL2_IIMM, `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)

`CASE_OP("ADD",   17'b0000000_000_0110011, `ALU_ADD,  `ALUSEL1_SRC1, `ALUSEL2_SRC2, `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("SUB",   17'b0100000_000_0110011, `ALU_SUB,  `ALUSEL1_SRC1, `ALUSEL2_SRC2, `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("SLL",   17'b0000000_001_0110011, `ALU_SLL,  `ALUSEL1_SRC1, `ALUSEL2_SRC2, `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("SLT",   17'b0000000_010_0110011, `ALU_SLT,  `ALUSEL1_SRC1, `ALUSEL2_SRC2, `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("SLTU",  17'b0000000_011_0110011, `ALU_SLTU, `ALUSEL1_SRC1, `ALUSEL2_SRC2, `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("XOR",   17'b0000000_100_0110011, `ALU_XOR,  `ALUSEL1_SRC1, `ALUSEL2_SRC2, `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("SRL",   17'b0000000_101_0110011, `ALU_SRL,  `ALUSEL1_SRC1, `ALUSEL2_SRC2, `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("SRA",   17'b0100000_101_0110011, `ALU_SRA,  `ALUSEL1_SRC1, `ALUSEL2_SRC2, `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("OR",    17'b0000000_110_0110011, `ALU_OR,   `ALUSEL1_SRC1, `ALUSEL2_SRC2, `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)
`CASE_OP("AND",   17'b0000000_111_0110011, `ALU_AND,  `ALUSEL1_SRC1, `ALUSEL2_SRC2, `WBSEL_ALURES, 1'b1, `CMP_X,    1'b0, 1'b0, 1'b0, 4'b0000)


`ifndef CMPOP
`define CMPOP

parameter [2:0] BEQ  = 0;
parameter [2:0] BNE  = 1;
parameter [2:0] BLT  = 2;
parameter [2:0] BGE  = 3;
parameter [2:0] BLTU = 4;
parameter [2:0] BGEU = 5;

`endif // CMPOP


`ifndef LSU
`define LSU

`define LSUOP_WIDTH 3
`define LSU_X      `LSUOP_WIDTH'dX
`define LSU_BYTE   `LSUOP_WIDTH'd0
`define LSU_HALF   `LSUOP_WIDTH'd1
`define LSU_WORD   `LSUOP_WIDTH'd2
`define LSU_U_BYTE `LSUOP_WIDTH'd3
`define LSU_U_HALF `LSUOP_WIDTH'd4

`endif // LSU


`ifndef OPCODE
`define OPCODE

parameter [3:0] ADD = 1;
parameter [3:0] SUB = 2;
parameter [3:0] SLL = 3;
parameter [3:0] SLT = 4;
parameter [3:0] SLTU= 5;
parameter [3:0] XOR = 6;
parameter [3:0] SRL = 7;
parameter [3:0] SRA = 8;
parameter [3:0] OR  = 9;
parameter [3:0] AND = 10;

`endif
